
/*
	reader of regFile,
	choose the right register output from 32 registers	
*/
/*
module regFileReader(input [4:0] ctrlReadReg,
							input [31:0] registerStates [31:0],
							output [31:0] selectedStates);
							
	// WRITE ME
	
	// YOU SHOULD USE THE triStateBuffer given
							

endmodule
*/